** Spice Models of Vishay 1 Mbd high speed optocouplers **
** Copyright VISHAY, Inc. 2010 All Rights Reserved.
**-- SFH6343T--**
* Same as 6N136  , w/o base
* Symbol Pin -> Model Node
*    A           1
*    K           2
*    E           3
*    C           4 
*    VCC         5 
.subckt SFH6343 A K GND C VCC
x1 A K GND C QB VCC 6N136
.ends SFH6343
*$
.SUBCKT 6N136  DA DK QE QC QB  VCC
DIN DA 9 DT8811VB
VT 9 DK 0
CIO DA QC 0.6e-12
QOUT QC QB QE QF290D
RFX QB QE 1e6
Hd T1 0 VT 800	;I-V
Rdly1 T1 T2 0.1
Cdly1 T2 0 1P
Gdly1 VCC QB VALUE {-2E-7 + 5e-6*V(T2) -1.7e-8*V(T2)*V(T2)}
.MODEL DT8811VB D 
+ IS=4.5E-18 N=1.40 RS=3.8
+ BV=3.000e+000 IBV=0.5e-006  XTI=4
+ EG=1.52436 CJO=18E-12 VJ=0.75 M=0.5 FC=0.5
.MODEL QF290D NPN 
+ IS=2.691e-016 NF=1.000e+000 ISE=6.586e-018
+ NE = 1.082e+000 BF = 176 BR = 1.000e+000
+ IKF = 7.300e-003 VAF = 1.000e+002 VAR = 2.800e+002
+ EG = 1.110e+000 XTI = 1.068e+000 XTB = 0.000e+000
+ RC = -1e+000 RB = 2.500e+001 RE = 40
+ CJE = 2.500e-012 MJE = 1.740e-001 VJE = 1.250e-001
+ CJC = 7.24e-012 MJC = 2.573e-001 VJC = 1.100e-001
.ENDS 6N136
