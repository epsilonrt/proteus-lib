*---------- DMG2305UX Spice Model ----------
.SUBCKT DMG2305UX 10 20 30 
*     TERMINALS:  D  G  S
M1 1 2 3 3 PMOS L = 1E-006 W = 1E-006 
RD 10 1 0.02969 
RS 30 3 0.001 
RG 20 2 15.2 
CGS 2 3 7.613E-010 
EGD 12 30 2 1 1 
VFB 14 30 0 
FFB 2 1 VFB 1 
CGD 13 14 1.28E-009 
R1 13 30 1 
D1 13 12 DLIM 
DDG 14 15 DCGD 
R2 12 15 1 
D2 30 15 DLIM 
DSD 10 3 DSUB 
.MODEL PMOS PMOS LEVEL = 3 U0 = 400 VMAX = 1E+006 ETA = 0.001 
+ TOX = 6E-008 NSUB = 1E+016 KP = 26.49 KAPPA = 65.74 VTO = -0.8201 
.MODEL DCGD D CJO = 5.79E-010 VJ = 0.2973 M = 0.5774 
.MODEL DSUB D IS = 3.162E-009 N = 1.241 RS = 0.08353 BV = 1E+006 CJO = 5.653E-011 VJ = 0.008286 M = 0.1128 
.MODEL DLIM D IS = 0.0001 
.ENDS
*Diodes DMG2305UX Spice Model v1.0 Last Revised 2013/10/22