*SRC=MMBT3904;DI_MMBT3904;BJTs NPN; Si; 40.0V 0.200A 347MHz Diodes Inc. NPN Transistor
.MODEL DI_MMBT3904 NPN (IS=48.3f NF=1.00 BF=410 VAF=114
+ IKF=0.121 ISE=13.1p NE=2.00 BR=4.00 NR=1.00
+ VAR=24.0 IKR=0.300 RE=2.63 RB=10.5 RC=1.05
+ XTB=1.5 CJE=9.67p VJE=1.10 MJE=0.500 CJC=8.70p VJC=0.300
+ MJC=0.300 TF=440p TR=74.7n EG=1.12 )