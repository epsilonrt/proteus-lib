*$
* Model: PS2715
*
* This SPICE model is intended to simulate the device behavior at Ta=25C within
* the maximum ratings as called out in the data sheet.
*
* Please note that the model can't duplicate exact device performance in the
* real world under all conditions and they can't replace the breadboarding 
* for final design verification.
*
* Note: CTR is modeled base on sample B in the data sheet. Please refer to the
* data sheet for details.
**********************************************************************************************
* A = PIN 1: diode anode
* K = PIN 2: diode cathode
* E = PIN 3: BJT emitter
* C = PIN 4: BJT collector
.SUBCKT PS2715 A K E C
D1 A D LED1
D2 F A LED2
Vsense1 D K 0
Vsense2 K F 0 
Hd1  J 0 Vsense1 1
Hd2  R J Vsense2 1
Rd   R T 100k
Cd   T 0 20p
Gctr C B TABLE
+ {If(V(T)<=5m,
+ ((-12780000000*PWR(V(T),5)+168500000*PWR(V(T),4)-
+ 850300*PWR(V(T),3)+2130*PWR(V(T),2)+0.9866*V(T)-0.0001351)*0.96/550),
+ ((886000*PWR(V(T),5)-148900*PWR(V(T),4)+
+ 9854*PWR(V(T),3)-315.9*PWR(V(T),2)+4.956*V(T)-0.001089)*0.98/550))}
+ (0,0) (0.1m, 0.1m) 
Q1 C B E detector
.model LED1 D IS=1p N=1.999644 RS=0 BV=6 IBV=10u
+ CJO=10p EG=1.424 TT=500n
.model LED2 D IS=1p N=1.999644 RS=0 BV=6 IBV=10u
+ CJO=10p EG=1.424 TT=500n
.model detector NPN IS=100p BF=550 NF=1.3 BR=50 TF=1n TR=1.5n
+ CJE=7p CJC=13p VAF=100 ISS=0 CJS=1p
.ends
*$
