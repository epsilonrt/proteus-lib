*
*DIODES_INC_SPICE_MODEL
*ORIGIN=DZSL_DPG_GM
*SIMULATOR=PSPICE
*DATE=10FEB2011
*VERSION=2
*PIN_ORDER         
* 1=C1    6=E1
* 2=B1    5=E2
* 3=B2    4=C2
*
.SUBCKT DMMT5401 1 2 3 4 5 6
Q1 1 2 6 Mod1
Q2 4 3 5 Mod1
*
.MODEL Mod1  PNP IS=6E-14 NF=1 BF=130 VAF=360 ISE=6E-14
+ NE=1.5 NR=1 BR=6.5 VAR=37 ISC=8E-12 NC=1.35 RC=0.08 RB=1 RE=0.25
+ CJC=13E-12 MJC=0.46  VJC=0.7 CJE=63E-12 MJE=0.41 VJE=0.9 
+ TF=6.7E-10 TR=1.03E-6 XTB=1.5 QUASIMOD=1 RCO=14 GAMMA=1.5E-8
.ENDS
*
*$