*ZETEX FZT600 Spice Model v1.0 Last Revised 23/12/04
*
.SUBCKT FZT600 1 2 3
*               C B E
Q1 1 2 4 SUB600
Q2 1 4 3 SUB600 2.74
*
.MODEL SUB600 NPN IS=8.354E-14 BF=70 VAF=18.3 IKF=0.25 ISE=2E-13
+NE=1.45 BR=2 VAR=6.5 NR=1 IKR=0.2 ISC=6.138E-13 NC=1.46 RB=0.5 RE=0.25
+RC=0.3 CJE=83.7E-12 VJE=0.6868 MJE=0.3362 CJC=8.6E-12 VJC=0.3679
+MJC=0.3607 TF=1E-9 TR=1800E-9
.ENDS FZT600
*
*$
*
