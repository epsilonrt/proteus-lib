** Spice3 of Vishay 1 Mbd high speed optocouplers **
** for parts: 6N136, 6N1136, SFH6136, SFH6316T, SFH6343T **
** Copyright VISHAY, Inc. 2010 All Rights Reserved.
* Symbol Pin -> Model Node
*    A           1
*    K           2
*    E           3
*    C           4
*    B           5 
*    VCC         6 
.SUBCKT 6N136 DA DK QE QC QB  VCC
DIN DA 9 DT8811VB
VT 9 DK 0
CIO DA QC 0.6e-12
QOUT QC QB QE QF290D
RFX QB QE 1e6
Hd T1 0 VT 800	;I-V
Rdly1 T1 T2 0.1
Cdly1 T2 0 1P
Gdly1 VCC QB VALUE {-2E-7 + 5e-6*V(T2) -1.7e-8*V(T2)*V(T2)}

.MODEL DT8811VB D 
+ IS=4.5E-18 N=1.40 RS=3.8
+ BV=3.000e+000 IBV=0.5e-006  XTI=4
+ EG=1.52436 CJO=18E-12 VJ=0.75 M=0.5 FC=0.5
.MODEL QF290D NPN 
+ IS=2.691e-016 NF=1.000e+000 ISE=6.586e-018
+ NE = 1.082e+000 BF = 176 BR = 1.000e+000
+ IKF = 7.300e-003 VAF = 1.000e+002 VAR = 2.800e+002
+ EG = 1.110e+000 XTI = 1.068e+000 XTB = 0.000e+000
+ RC = -1e+000 RB = 2.500e+001 RE = 40
+ CJE = 2.500e-012 MJE = 1.740e-001 VJE = 1.250e-001
+ CJC = 7.24e-012 MJC = 2.573e-001 VJC = 1.100e-001
.ENDS 6N136

**==================================================================*
* Note:                                                             *
* Altough models can be a useful tool in evaluating device          *
* performance, they cannot model exact device performance           *
* under all conditions, nor are they intended to replace            *
* breadboarding for final verification!                             *
*                                                                   *
* Models provided by VISHAY Semiconductors GmbH are not             *
* as fully representing all of the specifications and operating     *
* characteristics of the semiconductor product to which the         *
* model relates.                                                    *
* The models describe the characteristics of typical devices.       *
* In all cases, the current data sheet information for a given      *
* device is the final design guideline and the only actual          *
* performance specification.                                        *
* VISHAY Semiconductors does not assume any liability arising       *
* from the model use. VISHAY Semiconductors reserves the right to   *
* change models without prior notice.				        *
**==================================================================*
